module main

import peass2v

fn main() {
	peass2v.main_entry()
}